`timescale 1ns / 1ps

module MISR(CLK,RST,bist_end,e0,e1,e2,hf);
input CLK,RST,bist_end,e0,e1,e2;
reg h0,h1,h2,h3,h4,h5,h6,h7,h8,h9,h10,h11,h12,h13,h14,h15,h16,h17,h18,h19,h20 ;
output reg [20:0] hf;

always @(posedge CLK)
begin
    if (RST == 0)
    begin
    
        if (bist_end == 0) 
        begin
        h0 <= h1;
        h1 <= h2;
        h2 <= h3;
        h3 <= h4;
        h4 <= h5;
        h5 <= h6;
        h6 <= h7;
        h7 <= h8;
        h8 <= h9;
        h9 <= h10;
        h10 <= h11;
        h11 <= h12;
        h12 <= h13;
        h13 <= h14;
        h14 <= h15;
        h15 <= h16; 
        h16 <= h17;
        h17 <= h18;    
        h18 <= (e2 ^ h17);
        h19 <= (e1 ^ h18);
        h20 <= (e0 ^ (h19 ^ (h18 ^ (h17 ^ (h16 ^ (h15 ^ (h14 ^ (h13 ^ (h12 ^ (h11 ^ (h10 ^ (h9 ^ (h8 ^(h7 ^
                 (h6 ^(h5 ^(h4 ^(h3 ^ (h2 ^( h1 ^ h0 )))))))))))))))))))); 

//    h0 <= !(e2 || h1);
//    h1 <= !(e1 || h0); 
//    h2 <= !(e0 || !(h2 || !(h1||h0))); 
//    h3 <= !(h2 || h1);
//    h4 <= !(h3 || h2);
//    h5 <= !(h4 || h3);
//    h6 <= !(h5 || h4);
//    h7 <= !(h6 || h5);
//    h8 <= !(h7 || h6);
//    h9 <= !(h8 || h7); 
//    h10 <= !(h9 || h10);
//    h11 <= !(h10 || h9);
//    h12 <= !(h11 || h10);
//    h13 <= !(h12 || h11);
//    h14 <= !(h13 || h12);
//    h15 <= !(h14 || h11); 
//    h16 <= !(h15 || h12);
//    h17 <= !(h16 || h13);
//    h18 <= !(h17 || h14);
//    h19 <= !(h18 || h15);
//    h20 <= !(h19 || h16);
    hf <= {h0,h1,h2,h3,h4,h5,h6,h7,h8,h9,h10,h11,h12,h13,h14,h15,h16,h17,h18,h19,h20};
    end
    else
    h0 <= 1;
        h1 <= 1;
        h2 <= 1;
        h3 <= 1;
        h4 <= 1;
        h5 <= 1;
        h6 <= 1;
        h7 <= 1;
        h8 <= 1;
        h9 <= 1;
        h10 <= 1;
        h11 <= 1;
        h12 <= 1;
        h13 <= 1;
        h14 <= 1;
        h15 <= 1; 
        h16 <= 1;
        h17 <= 1;    
        h18 <= 1;
        h19 <= 1;
        h20 <= 1; 
        end
end
endmodule
